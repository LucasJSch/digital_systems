library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cordic_rotator is
end;

architecture cordic_rotator_arch of cordic_rotator is
end;